
module CPU(reset, clk);
	input reset, clk;
	
    //--------------Your code below-----------------------

    //...
        
    //--------------Your code above-----------------------

endmodule
	